module my_and(x1, x2, z);

input x1, x2;
output z;

    and a(z, x1, x2);

endmodule
